library verilog;
use verilog.vl_types.all;
entity HA_vlg_vec_tst is
end HA_vlg_vec_tst;
