library verilog;
use verilog.vl_types.all;
entity AccumulatorFINAL_vlg_vec_tst is
end AccumulatorFINAL_vlg_vec_tst;
