library verilog;
use verilog.vl_types.all;
entity ADDER_8_4_bits_vlg_vec_tst is
end ADDER_8_4_bits_vlg_vec_tst;
