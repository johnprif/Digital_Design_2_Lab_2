library verilog;
use verilog.vl_types.all;
entity FA_vlg_vec_tst is
end FA_vlg_vec_tst;
