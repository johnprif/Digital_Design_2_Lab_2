library verilog;
use verilog.vl_types.all;
entity AccumulatorOLD_vlg_vec_tst is
end AccumulatorOLD_vlg_vec_tst;
