library verilog;
use verilog.vl_types.all;
entity AccumulatorFINAL is
    port(
        Acc             : out    vl_logic_vector(7 downto 0);
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        ADD_SUB         : in     vl_logic;
        I               : in     vl_logic_vector(3 downto 0);
        Hex6            : out    vl_logic_vector(6 downto 0);
        Hex7            : out    vl_logic_vector(6 downto 0)
    );
end AccumulatorFINAL;
